module wallace_tree_reduction(a, b, r1, r2);
	input logic [5:0] a, b;
	output logic [11:0] r1, r2;
	// start your code here
endmodule
