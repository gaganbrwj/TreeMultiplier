module wallace_tree_reduction(a, b, r1, r2);
	input logic [4:0] a, b;
	output logic [9:0] r1, r2;
	// start your code here
endmodule
